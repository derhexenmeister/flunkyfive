//////////////////////////////////////////////////////////////////////
//
//////////////////////////////////////////////////////////////////////
`include "timescale.vh"
`include "ff_bfm_defines.vh"

module ff_utilities();
endmodule
