`timescale 1ns/100ps

// Use this to delay signals after a rising clock edge in simulation
// 
`ifndef D
    `define D   #1
`endif
